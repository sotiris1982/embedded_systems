interface clk_rstn_if;
	logic clk_i;
	logic rstn_i;
	
	
	
endinterface : clk_rstn_if